`ifndef BCD_ALU_OP_CODES_VH
`define BCD_ALU_OP_CODES_VH

`define BCD_ALU_OP_CODE_WIDTH 2

`define BCD_ALU_OP_SHL 2'h0
`define BCD_ALU_OP_SHR 2'h1
`define BCD_ALU_OP_ADD 2'h2
`define BCD_ALU_OP_CMP 2'h3

`endif
