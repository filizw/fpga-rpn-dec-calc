`ifndef BCDU_FLAGS_VH
`define BCDU_FLAGS_VH

`define BCDU_NUM_FLAGS 5

`define BCDU_ZF 0
`define BCDU_TF 1
`define BCDU_CF 2
`define BCDU_GF 3
`define BCDU_EF 4

`endif
