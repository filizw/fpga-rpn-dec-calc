`ifndef DAU_SYMBOLS_VH
`define DAU_SYMBOLS_VH

`define DAU_SYM_WIDTH 5

`define DAU_SYM_INVALID 5'h00

`define DAU_SYM_0 5'h10
`define DAU_SYM_1 5'h11
`define DAU_SYM_2 5'h12
`define DAU_SYM_3 5'h13
`define DAU_SYM_4 5'h14
`define DAU_SYM_5 5'h15
`define DAU_SYM_6 5'h16
`define DAU_SYM_7 5'h17
`define DAU_SYM_8 5'h18
`define DAU_SYM_9 5'h19

`define DAU_SYM_COMMA 5'h1C

`define DAU_SYM_PLUS  5'h1B
`define DAU_SYM_MINUS 5'h1D

`define DAU_SYM_MUL 5'h1A
`define DAU_SYM_DIV 5'h1F

`define DAU_SYM_SEPARATOR 5'h02
`define DAU_SYM_RESULT    5'h0D
`define DAU_SYM_NEW_LINE  5'h0A
`define DAU_SYM_RESET     5'h07

`endif
