`ifndef BCDU_OP_CODES_VH
`define BCDU_OP_CODES_VH

`define BCDU_OP_CODE_WIDTH 4

`define BCDU_OP_NOP 4'h0
`define BCDU_OP_SHL 4'h1
`define BCDU_OP_SHR 4'h2
`define BCDU_OP_ADD 4'h3
`define BCDU_OP_SUB 4'h4
`define BCDU_OP_CMP 4'h5
`define BCDU_OP_CLR 4'h6
`define BCDU_OP_MOV 4'h7
`define BCDU_OP_ACA 4'h8
`define BCDU_OP_ACS 4'h9

`endif
